module main

fn test_dummy() {
	assert true
}
